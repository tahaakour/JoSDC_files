// Code your design here
module and32(in1 , in2 , out);
  
  input [31:0] in1,in2;
  output [31:0] out;
  
  wire [31:0] in1_w, in2_w;
  
  assign in1_w = in1;
  assign in2_w = in2;
  
  
  assign out = in1 & in2;
  
endmodule

  